-------------------------------------------------------------------------------
--
-- Title       : SixBitProcessorWithMultiplier
-- Design      : SixBitProcessor
-- Author      : Alireza
-- Company     : AC
--
-------------------------------------------------------------------------------
--
-- File        : C:\Users\zephyrus\Desktop\CoDes_Project_Changiziyan_Alireza_Salehi_Sadra\CoDesProject\SixBitProcessor\src\SixBitProcessorWithMultiplier.vhd
-- Generated   : Thu Jul  4 15:32:03 2024
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {SixBitProcessorWithMultiplier} architecture {SixBitProcessorWithMultiplier}}



entity SixBitProcessorWithMultiplier is
end SixBitProcessorWithMultiplier;

--}} End of automatically maintained section

architecture SixBitProcessorWithMultiplier of SixBitProcessorWithMultiplier is
begin

	 -- enter your statements here --

end SixBitProcessorWithMultiplier;
